`define EXAMPLE_CONSTANT 10
